
module nios_td3 (
	clk_clk,
	reset_reset_n,
	pio_0_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	pio_0_export;
endmodule
