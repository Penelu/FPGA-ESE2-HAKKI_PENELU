// nios_td3_tb.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module nios_td3_tb (
	);

	wire    nios_td3_inst_clk_bfm_clk_clk;       // nios_td3_inst_clk_bfm:clk -> [nios_td3_inst:clk_clk, nios_td3_inst_reset_bfm:clk]
	wire    nios_td3_inst_reset_bfm_reset_reset; // nios_td3_inst_reset_bfm:reset -> nios_td3_inst:reset_reset_n

	nios_td3 nios_td3_inst (
		.clk_clk       (nios_td3_inst_clk_bfm_clk_clk),       //   clk.clk
		.pio_0_export  (),                                    // pio_0.export
		.reset_reset_n (nios_td3_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_td3_inst_clk_bfm (
		.clk (nios_td3_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nios_td3_inst_reset_bfm (
		.reset (nios_td3_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nios_td3_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
